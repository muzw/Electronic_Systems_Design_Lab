-- FPGA_EXP4_mzw @ PB20051061

